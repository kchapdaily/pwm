----------------------------------------------------------------------------------
-- Company: 
-- Engineer: KEVIN CHAPMAN
-- 
-- Create Date:    21:13:23 05/16/2013 
-- Design Name: 
-- Module Name:    top_level_pwm - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity top_level_pwm is
end top_level_pwm;

architecture Behavioral of top_level_pwm is

begin


end Behavioral;

